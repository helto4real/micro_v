module binding

import lib.comp.types

[heap]
pub struct VariableSymbol {
pub:
	name   string
	typ    types.Type
	is_mut bool
}

pub fn (vs &VariableSymbol) str() string {
	mut_str := if vs.is_mut {'mut '} else {''}
	return 'VariableSymbol $mut_str <$vs.name> ($vs.typ)'
}

pub fn new_variable_symbol(name string, typ types.Type, is_mut bool) &VariableSymbol {
	return &VariableSymbol {
		name: name
		typ: typ
		is_mut: is_mut
	}
}