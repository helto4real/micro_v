module v
import parser
import token

pub struct Compiler {

}

pub fn new_compiler(args Arg) &Compiler {
	return &Compiler {}
}