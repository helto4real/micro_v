// bidning module binds to the syntax tree and handle checks
module binding

import lib.comp.ast
import lib.comp.util

[heap]
pub struct Binder {
pub mut:
	scope &BoundScope
	log   &util.Diagnostics // errors when parsing
}

pub fn new_binder(parent &BoundScope) &Binder {
	return &Binder{
		scope: new_bound_scope(parent)
		log: util.new_diagonistics()
	}
}

pub fn bind_global_scope(previous &BoundGlobalScope, comp_node &ast.ComplationSyntax) &BoundGlobalScope {
	parent_scope := create_parent_scope(previous)
	mut binder := new_binder(parent_scope)
	stmt := binder.bind_stmt(comp_node.stmt)
	vars := binder.scope.vars()
	mut diagnostics := binder.log.all
	if previous != 0 && previous.log.all.len > 0 {
		diagnostics.prepend(previous.log.all)
	}
	return new_bound_global_scope(previous, binder.log, vars, stmt)
}

fn create_parent_scope(previous &BoundGlobalScope) &BoundScope {
	mut stack := new_bound_global_scope_stack()
	mut prev := previous

	for prev != 0 {
		stack.push(prev)
		prev = prev.previous
	}
	mut parent := &BoundScope(0)

	for !stack.is_empty() {
		prev = stack.pop() or { &BoundGlobalScope(0) }
		if prev == 0 {
			panic('unexpected return from stack')
		}
		mut scope := new_bound_scope(parent)
		for var in prev.vars {
			scope.try_declare(var)
		}
		parent = scope
	}

	return parent
}

pub fn (mut b Binder) bind_stmt(stmt ast.StatementSyntax) BoundStmt {
	match stmt {
		ast.BlockStatementSyntax { return b.bind_block_stmt(stmt) }
		ast.ExpressionStatementSyntax { return b.bind_expr_stmt(stmt) }
		ast.VarDeclStmtSyntax { return b.bind_var_decl_stmt(stmt) }
		ast.IfStmtSyntax { return b.bind_if_stmt(stmt) }
	}
}
pub fn (mut b Binder) bind_if_stmt(if_stmt ast.IfStmtSyntax) BoundStmt {
	return BoundStmt{}
}

pub fn (mut b Binder) bind_block_stmt(block_stmt ast.BlockStatementSyntax) BoundStmt {
	b.scope = new_bound_scope(b.scope)
	mut stmts := []BoundStmt{}
	for i, _ in block_stmt.statements {
		stmts << b.bind_stmt(block_stmt.statements[i])
	}
	b.scope = b.scope.parent
	return new_bound_block_stmt(stmts)
}

pub fn (mut b Binder) bind_expr_stmt(expr_stmt ast.ExpressionStatementSyntax) BoundStmt {
	expr := b.bind_expr(expr_stmt.expr)
	return new_bound_expr_stmt(expr)
}

pub fn (mut b Binder) bind_expr(expr ast.ExpressionSyntax) BoundExpr {
	match expr {
		ast.LiteralExpr { return b.bind_literal_expr(expr) }
		ast.UnaryExpr { return b.bind_unary_expr(expr) }
		ast.BinaryExpr { return b.bind_binary_expr(expr) }
		ast.ParaExpr { return b.bind_para_expr(expr) }
		ast.NameExpr { return b.bind_name_expr(expr) }
		ast.AssignExpr { return b.bind_assign_expr(expr) }
		else { panic('unexpected bound expression $expr') }
	}
}

pub fn (mut b Binder) bind_var_decl_stmt(syntax ast.VarDeclStmtSyntax) BoundStmt {
	name := syntax.ident.lit
	bound_expr := b.bind_expr(syntax.expr)

	var := new_variable_symbol(name, bound_expr.typ(), syntax.is_mut)
	res := b.scope.try_declare(var)
	if res == false {
		b.log.error_name_already_defined(name, syntax.ident.pos)
	}
	return new_var_decl_stmt(var, bound_expr, syntax.is_mut)
}

fn (mut b Binder) bind_assign_expr(syntax ast.AssignExpr) BoundExpr {
	name := syntax.ident.lit
	bound_expr := b.bind_expr(syntax.expr)

	// check is varable exist in scope
	mut var := b.scope.lookup(name) or {
		// var have to be declared with := to be able to set a value
		b.log.error_var_not_exists(name, syntax.ident.pos)
		return bound_expr
	}

	if !var.is_mut {
		// trying to assign a nom a mutable var
		b.log.error_assign_non_mutable_variable(name, syntax.eq_tok.pos)
	}

	if bound_expr.typ() != var.typ {
		b.log.error_cannot_convert_variable_type(bound_expr.typ_str(), var.typ.typ_str(),
			syntax.expr.pos())
		return bound_expr
	}
	return new_bound_assign_expr(var, bound_expr)
}

fn (mut b Binder) bind_para_expr(syntax ast.ParaExpr) BoundExpr {
	return b.bind_expr(syntax.expr)
}

fn (mut b Binder) bind_name_expr(syntax ast.NameExpr) BoundExpr {
	name := syntax.ident_tok.lit
	variable := b.scope.lookup(name) or {
		b.log.error_var_not_exists(name, syntax.ident_tok.pos)
		return new_bound_literal_expr(0)
	}
	return new_bound_variable_expr(variable)
}

fn (mut b Binder) bind_literal_expr(syntax ast.LiteralExpr) BoundExpr {
	val := syntax.val
	return new_bound_literal_expr(val)
}
