module util

pub struct Pos {
pub:
	pos int // position in textfile
	ln  int // line number
	col int // column of line
}