fn main() {
	println('hello world!')
}

module test
main()
