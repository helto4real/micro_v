module args

pub struct Args {
}
