module my_mod 

fn a_cool_module(i int) int {
	return i
}