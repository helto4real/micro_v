module util

pub struct Message {
pub:
	pos  Pos    // position of error
	text string // error text
}