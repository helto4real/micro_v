module parser

pub struct Parser {
	
}