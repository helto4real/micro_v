module comp

pub struct Args {
}
